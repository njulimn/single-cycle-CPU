module I_mm_read(I_mem_addr,IR);


input [31:0]  	 	I_mem_addr;
output  reg [31:0]   		IR;


reg  [7:0] inst[63:0];
	
  initial
	begin
		{inst[3],inst[2],inst[1],inst[0]} =    	32'b000000_00001_00010_00011000_00100000;       	 //add   R3 = R1+R2
		{inst[7],inst[6],inst[5],inst[4]} = 		32'b001000_00100_00111_00000000_10000000;     		 //addi  R7 = R4+128
		{inst[11],inst[10],inst[9],inst[8]} = 		32'b001001_00100_01000_00000000_10000000;     		 //addiu R8 = R4+128
		{inst[15],inst[14],inst[13],inst[12]} = 	32'b000000_00001_00010_01001000_00100010;   		 	 //sub   R9 = R1-R2
		
		{inst[19],inst[18],inst[17],inst[16]} = 	32'b000000_00001_00010_01010000_00100011;     	 	 //subu  R10 = R1-R2
		{inst[23],inst[22],inst[21],inst[20]} = 	32'b011111_00000_00001_11000_00010_100000;   		 //seb   R1 R24
		{inst[27],inst[26],inst[25],inst[24]} = 	32'b001111_00000_10000_0101010101010101;   	 	 	 //lui  R16    0101010101010101 
		{inst[31],inst[30],inst[29],inst[28]} = 	32'b001110_00001_01100_0101010101010101;   		  	 //xori  R12 = R1^0101010101010101
		
		{inst[35],inst[34],inst[33],inst[32]} = 	32'b011100_00001_00000_01101_00000_100001;   		 //clo   R13 = clo R1
		{inst[39],inst[38],inst[37],inst[36]} = 	32'b011100_00010_00000_01110_00000_100000;   	    //clz   R14 = clz R2
		{inst[43],inst[42],inst[41],inst[40]} = 	32'b000000_00101_00100_10000_00000_000111;   		 //SRAV  R16 R4>>5=R32;
		{inst[47],inst[46],inst[45],inst[44]} = 	32'b000000_0000_1_00101_10000_00100_000010;   		 //rotr  R16 R5>>4(shmat);
		
		{inst[51],inst[50],inst[49],inst[48]} = 	32'b000000_00001_00010_10000_00000_101011;   		 //sltu  R16 = R1<R2
		{inst[55],inst[54],inst[53],inst[52]} = 	32'b001010_00001_10001_1111111111111111;   		    //slti  R17 = R1<32767   
		{inst[59],inst[58],inst[57],inst[56]} = 	32'b000010_00000000000000000000001111;   		       //j      60
		{inst[63],inst[62],inst[61],inst[60]} = 	32'b000001_00001_11111_0000000000000001;   			 //bgez  R1 OFFSET 1      
		
	end


always @ (*)
	begin
		IR[7:0] 		= inst[I_mem_addr];
		IR[15:8] 	= inst[I_mem_addr+1];
		IR[23:16] 	= inst[I_mem_addr+2];
		IR[31:24] 	= inst[I_mem_addr+3];
	end

endmodule


